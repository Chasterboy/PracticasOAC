library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity concatenador_datos is
	Port(entradaA : in STD_LOGIC_VECTOR(2 downto 0); --Entrada
			entradaB: in STD_LOGIC_VECTOR(2 downto 0); --Edo siguiente
			salida : out STD_LOGIC_VECTOR(5 downto 0));
end concatenador_datos;

architecture Behavioral of concatenador_datos is
begin
		process(entradaA, entradaB)
		begin
			salida <= entradaB & entradaA; --Liga & Entradas
		end process;
end Behavioral;
		