library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is
Port ( 
	dir : in STD_LOGIC_VECTOR (11 downto 0);
	data : out STD_LOGIC_VECTOR (97 downto 0));
end memory;

architecture Behavioral of memory is

begin
	process(dir)
	begin
	
		-- DATA FORMAT
		-- |    PRUEBA    |VF| Ins |                LIGA                 |
		--  P4 P3 P2 P1 P0 VF I1 I0 L11 L10 L9 L8 L7 L6 L5 L4 L3 L2 L1 L0 nCRI EB1 EB0 nWB EA1 EA0 nWA selbus UPA9 UPA8 UPA7 UPA6 UPA5 UPA4 UPA3 UPA2 UPA1 UPA0 nOEUPA nDUPA selmux nEX2 nEX1 nEX0 X2 X1 X0 EnaY nERA2 nERA1 nERA0 RA2 RA1 RA0 nEAP2 nEAP1 nEAP0 AP2 AP1 AP0 nEPC2 nEPC1 nEPC0 PC2 PC1 PC0 nCBD nAS nRW BD DINT HINT SET_IRQ SET_XIRQ B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 CC CN CV CZ CI CH CX CS nHB ACCSEC

		-- Cadena por default: "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010"
		
		--if(dir=    X"000") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";
		--elsif(dir= X"001") then data <= "00000" & "0" & "00" & "000000000000" & "00000000000000000000000000000000000000000000000000000000000000000000000000"; 
												  
		--Fetch										  
		if(dir=    X"000") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"001") then data <= "00000000000000000000000100100000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"002") then data <= "00000010000000000000100100100000000000110111000011100011100011100011111110000000000000000000000010";

		--LDAA (INM)
		elsif(dir= X"860") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"861") then data <= "00000000000000000000100101000000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"862") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"863") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--LDAB (INM)
		elsif(dir= X"C60") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"C61") then data <= "00000000000000000000101000100000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"C62") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000100101000111000010";
		elsif(dir= X"C63") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--ABA (INH)
		elsif(dir= X"1B0") then data <= "00000000000000000000111111100000000001111111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"1B1") then data <= "01111111000000000000100101000000000000000111000011100011100011100011111110000000000000001111010010";
		elsif(dir= X"1B2") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--JMP (EXT)
		elsif(dir= X"7E0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7E1") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"7E2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7E3") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"7E4") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111110000000000000000000000010";
		elsif(dir= X"7E5") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--CMP (INH)
		elsif(dir= X"1A0") then data <= "00000000000000000000111111100000100001111111000011100011100011100011111110000000000000000000000011";
		elsif(dir= X"1A1") then data <= "01111111000000000000100100100000000000000111000011100011100011100011111110000000000000001111010010";
		elsif(dir= X"1A2") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--JB (EXT)
		elsif(dir= X"080") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"081") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"082") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"083") then data <= "10011001000010000101100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"084") then data <= "01111100000000000000100100100000000000110111000010000011100010010111111110000000000000000000000010";
		elsif(dir= X"085") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--JE (EXT)
		elsif(dir= X"7D0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7D1") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"7D2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7D3") then data <= "10010001011111010101100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"7D4") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111010000000000000000000000010";
		elsif(dir= X"7D5") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--Jc (EXT)
		elsif(dir= X"670") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"671") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"672") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"673") then data <= "10000001011001110101100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"674") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111010000000000000000000000010";
		elsif(dir= X"675") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--STAA (EXT)
		elsif(dir= X"A70") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"A71") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111010000000000000000000000010";
		elsif(dir= X"A72") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"A73") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"A74") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"A75") then data <= "00000000000000000000100101100000000000110111000011100011100011100011111000000000000000000000000010";
		elsif(dir= X"A76") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"A77") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--LDAA (EXT)
		elsif(dir= X"760") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"761") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111010000000000000000000000010";
		elsif(dir= X"762") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"763") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"764") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"765") then data <= "00000000000000000000100101000000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"766") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"767") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--LDAB (EXT)
		elsif(dir= X"B60") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"B61") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111010000000000000000000000010";
		elsif(dir= X"B62") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"B63") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"B64") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"B65") then data <= "00000000000000000000101000100000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"B66") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"B67") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--STAA (DIR)
		elsif(dir= X"A80") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"A81") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir= X"A82") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"A83") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"A84") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"A85") then data <= "00000000000000000000100101100000000000110111000011100011100011100011111000000000000000000000000010";
		elsif(dir= X"A86") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"A87") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--LDAA (DIR)
		elsif(dir= X"960") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"961") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir= X"962") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"963") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"964") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"965") then data <= "00000000000000000000100101000000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"966") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"967") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--LDAB (DIR)
		elsif(dir= X"D60") then data <= "00000000000000000000111100100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"D61") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir= X"D62") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"D63") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"D64") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"D65") then data <= "00000000000000000000101000100000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"D66") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"D67") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--STAA (IND)
		elsif(dir= X"A90") then data <= "00000000000000000000100100100000000000110111000011001101100011100001111110000000000000000000000000";
		elsif(dir= X"A91") then data <= "00000000000000000000100100100000110111110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"A92") then data <= "00000000000000000000100100100010000110111110000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"A93") then data <= "00000101101010011011100100100000000000000110011011100011100011100011111110000000000000001000000010";
		elsif(dir= X"A94") then data <= "00000000000000000000100100110010000111110101000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"A95") then data <= "00000000000000000000100100100000000000000101100011100011100011100011111110000000000000000000000010";
		elsif(dir= X"A96") then data <= "00000000000000000000100100100000000000110111100011000011100011100011111110000000000000011000000000";
		elsif(dir= X"A97") then data <= "00000000000000000000100100100000000000110011000011100011100011100001111110000000000000000000000010";
		elsif(dir= X"A98") then data <= "00000000000000000000100101100000000000110111000011100011100011100011111000000000000000000000000010";
		elsif(dir= X"A99") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"A9A") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"A9B") then data <= "11000001101010010101100100110010100111110101000011100011100011100011111110000000000000000000000010";
		
		--LDAA (IND)
		elsif(dir= X"A60") then data <= "00000000000000000000100100100000000000110111000011001111100001100001111110000000000000000000000000";
		elsif(dir= X"A61") then data <= "00000000000000000000100100100000110111110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"A62") then data <= "00000000000000000000100100100010000110111110000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"A63") then data <= "00000001101001101011100100100000000000000110011011100011100011100011111110000000000000001000000010";
		elsif(dir= X"A64") then data <= "00000000000000000000100100110010000111110111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"A65") then data <= "00000000000000000000100100100000000000000101100011100011100011100011111110000000000000000000000010";
		elsif(dir= X"A66") then data <= "00000000000000000000100100100000000000110111100011000011100011100011111110000000000000011000000000";
		elsif(dir= X"A67") then data <= "00000000000000000000100100100000000000110011000011100011100011100001111110000000000000000000000010";
		elsif(dir= X"A68") then data <= "00000000000000000000100101000000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"A69") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"A6A") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"A6B") then data <= "11000001101001100101100100110010100111110101000011100011100011100011111110000000000000000000000010";
		
		--LDAB (IND)
		elsif(dir= X"E60") then data <= "00000000000000000000100100100000000000110111000011001111100001100001111110000000000000000000000000";
		elsif(dir= X"E61") then data <= "00000000000000000000100100100000110111110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"E62") then data <= "00000000000000000000100100100010000110111110000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"E63") then data <= "00000101111001101011100100100000000000000110011011100011100011100011111110000000000000001000000010";
		elsif(dir= X"E64") then data <= "00000000000000000000100100110010000111110101000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"E65") then data <= "00000000000000000000100100100000000000000101100011100011100011100011111110000000000000000000000010";
		elsif(dir= X"E66") then data <= "00000000000000000000100100100000000000110111100011000011100011100011111110000000000000011000000000";
		elsif(dir= X"E67") then data <= "00000000000000000000100100100000000000110011000011100011100011100001111110000000000000000000000010";
		elsif(dir= X"E68") then data <= "00000000000000000000101000100000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"E69") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"E6A") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"E6B") then data <= "11000001111001100101100100110010100111110101000011100011100011100011111110000000000000000000000010";
		
	
		elsif(dir= X"200") then data <= "11000001000000000000100100100000000000110111000011100011100010010111011110000000000000000000000010";
		
		--else data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000000000000000000010"; -- Default
		else data <= "00000000000000000000100100100000000000110111000011100011100011100011111110000000000000000000000010";

		end if;
	end process;
end Behavioral;