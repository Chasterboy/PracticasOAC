LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY mux_entradas IS
    PORT (
        Sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        I0 : IN STD_LOGIC; --
        I1 : IN STD_LOGIC; --
        I2 : IN STD_LOGIC; --
        I3 : IN STD_LOGIC; --
        L : out STD_LOGIC 
    );
END mux_entradas;
ARCHITECTURE Behavioral OF mux_entradas IS
BEGIN
    PROCESS (Sel, I0, I1, I2, I3)
    BEGIN
        IF Sel = "00" THEN
            L <= I0;
        ELSIF Sel = "01" THEN
            L <= I1;
        ELSIF Sel = "10" THEN
            L <= I2;
        ELSIF Sel = "11" THEN
            L <= I3;
        END IF;
    END PROCESS;
END Behavioral;